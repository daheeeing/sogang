`timescale 1ns / 1ps

module bcd_adder_tb;
    reg [3:0] A, B;
    reg Cin;
    wire [7:0] S;
    wire [6:0] C;
    wire Cout, K;
    
bcd_adder u_bcd_adder(
    .A(A),
    .B(B),
    .Cin(Cin),
    .S(S),
    .C(C),
    .Cout(Cout),
    .K(K)
);

initial A = 4'D0;
initial B = 4'D0;
initial Cin = 1'b0;

always@(A or B or Cin)begin
A <= #10 A+4'D1;
B <= #20 A-4'D1;
Cin <= #30 ~Cin;
end

initial begin
    #1500
    $finish;
end
endmodule
